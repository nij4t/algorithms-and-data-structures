module main

fn main() {
	println('vello world!')
}